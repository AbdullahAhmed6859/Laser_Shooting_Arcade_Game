`timescale 1ns / 1ps

module clk_div (clk, clk_d);
    parameter div_value = 4999;
    input clk;
    output clk_d;
    reg clk_d;
    reg [19:0] count;
    initial begin
    clk_d = 1'b0; 
    count = 0;
    end
    always @(posedge clk) begin
        if (count == div_value) begin
        count <= 0; // reset count
        clk_d <= ~ clk_d;
        end else begin
        count <= count + 1; // count up
        end
    end
endmodule